`timescale 1 ns / 1 ps
module tb_lbp();
    

endmodule
